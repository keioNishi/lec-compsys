module ackor(input a0, a1, a2, a3, output ao);
	assign ao = a0 | a1 | a2 | a3;
endmodule
