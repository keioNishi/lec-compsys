`include "sw.vh"
module isbm(input [1:0] pout, output logic re, input empty,
	input [`PORT:0] reqi, output logic [`PORT:0] req, input ack, input clk, rst);
	typedef enum {INIT, AREQ, XFER} ISBMTYPE;
	ISBMTYPE state, nstate;
//
//
//
//
//
//
//
//
//
endmodule
