module test(a, b);
	output b;
	input a;
	assign b = a;
endmodule
